asearch.AND=OCH
asearch.AdvancedSearch=Avancerad sökning
asearch.All=Alla
asearch.AllDataProviders=Alla dataleverantörer
asearch.Between=Mellan
asearch.Contains=Innehåller
asearch.NOT=EJ
asearch.OR=ELLER
asearch.SearchIn=Sök i
asearch.Select=Välj
asearch.SelectDataProviders=Välj dataleverantör
cms.AddPageToAMenu=Lägg till sidan i en meny
cms.AddingImages=Lägg till bilder
cms.AreYouSureYouWantToDelete=Är du säker på att du vill ta bort denna sida och alla versioner av den? Detta kan inte ångras.
cms.AutoGeneratePageKey=Auto-generera sidnamn
cms.BeginByChoosingAnImage=<ul><li>Börja med att välja bild från din dator genom att trycka <span class="btn btn-success btn-mini"><i class="icon-plus icon-white"></i>Välj en bild</span></li><li>Du kan välja en eller fler bilder</li></ul>
cms.CreateANewPage=Skapa ny sida
cms.CreatingContentForTheHomePage=Att skapa en hemsida fungerar exakt likadant som att skapa en vanlig sida förutom följande: <ol><li><strong>Sidnnamnet</strong> måste vara: <em>hemsida</em></li><li>Sidan kan inte läggas till en meny</li></ol>
cms.CreatingHomepageContent=Skapa innehåll för hemsidan
cms.DeletePage=Ta bort sida
cms.FieldsExplained=Fältförklaring
cms.HelpWithUploadingImages=Hjälp att ladda upp bilder
cms.HelpWithWebsitePages=Hjälp med webbsidor
cms.Homepage=Hemsida
cms.ImagesCanBeAdded=Bilder kan läggas till på två sätt: <ol><li><strong>Ladda upp från en dator:</strong> detta kan du göra på <a href="/organizations/{0}/site/upload">Ladda upp bild</a> sidan. När bilden sparats kan den användas i din webbsida genom att klicka på <span class="mceIcon mceImage"></span> ikonen och välj din bild i <em>bildlistan</em></li><li><strong>Direkt från Internet:</strong> Klicka på <span class="mceIcon mceImage"></span> ikonen och skriv in webbadressen till bilden i </em>Bild URL</em> fältet
cms.InvalidKeyValue=Felaktig inmatning. Sidnamnet får bara vara med små bokstäver och mellan 3 och 35 tecken långt.
cms.ListPagesIn=Lista sidor i 
cms.MainMenu=Huvudmeny
cms.MakeThisContentAvailable=Om du kryssar i här gör du innehållet publikt
cms.NotPublished=Ej publicerad
cms.OnceUploaded=<p>När du har laddat upp, gå tillbaks till <a href="/organizations/{0}/site">sidlista</a> och redigera en sida eller skapa en <a href="/organizations/{0}/site/{1}/page/add">ny sida</a>. Klicka på <span class="mceIcon mceImage"></span> ikonen för att välja bild från <em>bildlistan</em>.</p>
cms.PageKey=Sidnamn
cms.PositionInTheMenu=Position i menyn
cms.Publish=Publicera
cms.Published=Publicerad
cms.ReadyForUse=Klar att använda
cms.SaveFiles=Spara filer
cms.SavePage=Spara sida
cms.SelectTheMenu=Välj menyn du vill att sidlänken ska visas i.
cms.SiteContentAdministrationRights=Administratörsrättigheter på sidinnehåll
cms.TheHubTheme=Hubtemat för denna sida.
cms.TheImagesAreThenAdded=<p>Bilderna är sedan tillagda och kan laddas upp till CultureHub.</p><ul><li>Klicka på <span class="btn btn-primary btn-mini"><i class="icon-upload icon-white"></i>Ladda upp</span> för att ladda upp alla bilder</li><li>Klicka på <span class="btn btn-primary btn-mini"><i class="icon-upload icon-white"></i>Ladda upp</span> på varje bild i listan för att ladda upp bilderna en och en</li></ul>
cms.TheLanguageOfThisPage=Språk för aktuell sida. Om språkväxling är aktivt (om du har flerspråksstöd i din Hub) bör du skapa en sida för varje språk.
cms.ThePositionOfYourPageLink=Positionen på sidlänken i vald meny. Ju högre nummer, ju längre till höger flyttar den.
cms.TitleMandatory=Titel måste finnas för sidnamnsgenerering.
cms.UniqueIdentifierForThePage=Unikt id för sidan. Detta id används som URL för sidan.
cms.UpdateHomepage=Uppdatera hemsidan
cms.UpdatePage=Uppdatera sidan
cms.UploadFile=Ladda upp filer
cms.UploadImage=Ladda upp bilder
cms.UsedInThePagesHTML=Används i sidans html <code>&lt;title&gt;&lt;/title&gt;</code> attribut, och om sidan är tillagd i menyn kommer detta med som länk i menyn.
cms.UsingTemplates=Använder mallar
cms.WebsitePages=Webbsidor
cms.WhenCreatingPageContent=När du skapar en sida går det snabbare om du använder en mall. Klicka på <span class="mceIcon mceTemplate"></span> ikonen så öppnas ett fönster där du kan granska och välja mallar
dataset.AreYouSureYouWantToRemoveThisDataset=Är du säker på att du vill radera datasetet?
dataset.BeginTypingADatasetName=Börja ange ett namn på datasetet
dataset.CancelProcessing=Avbryt bearbetningen
dataset.CannotAddDatasetWithId=Kan inte lägga till datasetet med id {0} till gruppen {0}
dataset.CreateADataset=Skapa ett dataset
dataset.CreateNewDatasetForUser=Skapa nytt dataset för användare {0}
dataset.DataSetWasNotFound=Dataset {0} hittades inte
dataset.Dataset=Dataset
dataset.DatasetCannotBeDeleted=Datasetet kan inte raderas just nu
dataset.DatasetCannotBeDisabled=Datasetet kan inte inaktiveras just nu
dataset.DatasetCannotBeEnabled=Datasetet kan inte aktiveras just nu
dataset.DatasetCannotBeProcessed=Datasetet kan inte bearbetas just nu
dataset.DatasetCannotBeReProcessed=Datasetet kan inte ombearbetas just nu
dataset.DatasetHashesCannotBeReset=Datasetets hashar kan inte återställas just nu
dataset.DatasetIndexingCannotBeCancelled=Datasetets indexering kan inte avbrytas just nu
dataset.DatasetInformation=Dataset Information
dataset.DatasetList=Dataset lista
dataset.DatasetWasNotFound=Dataset {0} hittades inte
dataset.Datasets=Dataset 
dataset.Disable=Inaktivera
dataset.Disabled=Inaktiverad
dataset.Enable=Aktivera
dataset.Enabled=Aktiverad
dataset.ErrorOccurredWhileProcessing=Det uppstod fel vid bearbetningen
dataset.FilterByName=Filtrera på namn
dataset.FilterByState=Filtrera på status
dataset.FindADataset=Find a dataset
dataset.Identifier=Identifierare
dataset.Incomplete=Ofullständig
dataset.ListOfDatasets=Lista över dataset
dataset.ListOfDatasetsForUser=Lista över dataset för användare {0}
dataset.Locked=Låst
dataset.LockedBy=Låst av:
dataset.NumberDatasets={0} Dataset(s)
dataset.NumberOfDatasets=Antal Dataset
dataset.ParsingAndStoring=Analysering och lagring av uppladdat data
dataset.Process=Bearbeta
dataset.Processing=Bearbetning
dataset.ProcessingCancelled=Bearbetning avbruten
dataset.QueuedForProcessing=I kö för bearbetning
dataset.ReProcess=Ombearbeta
dataset.ResetHashes=Återställ hashes
dataset.SaveDataset=Spara Dataset
dataset.TheQuotaOfAllowedDatasetsExceeded=Kvoten för antal tillåtna Dataset för denna organisation har överskridits
dataset.TheUniqueIdentifierOfThisDataset=Unikt id för detta Dataset
dataset.ThisDatasetIdentifierIsAlreadyInUse=Detta Dataset id används redan
dataset.Unlocked=Olåst
dataset.UpdateADataset=Uppdatera ett dataset
dataset.UpdateDatasetForUser=Uppdatera dataset för användare {0}
dataset.UploadedAndReady=Uppladdad och redo för bearbetning 
dataset.YouNeedToDisableTheDataset=Du måste inaktivera datasetet innan det kan raderas
hub.AFewWordsAboutYourself=Några ord om dig själv
hub.AboutYou=Om dig
hub.AccountSpace=Kontots utrymme
hub.Add=Lägg till
hub.AddANewMember=Lägg till en ny medlem genom att skriva användarnamnet i det tomma fältet ovanför och tryck ENTER.
hub.AddAnAdministrator=Lägg till en administratör genom att skriva användarnamnet i det tomma fältet ovanför och tryck ENTER.
hub.AddComment=Lägg till kommentar
hub.AddFiles=Lägg till filer...
hub.AddLabel=Lägg till etikett
hub.Administration=Administration
hub.AdministratorOptions=Administratörsalternativ
hub.AdministratorRights=Administratörsrättigheter
hub.Administrators=Administratörer
hub.All=Alla
hub.AlsoIncludeResultsWithoutImages=Ta även med poster utan bild
hub.AnEmailHasBeenSentToResetYourPassword=Ett e-postmeddelande har skickats till dig med en länk för att återställa lösenordet
hub.AreYouSureYouWantToDeleteThisGroup=Är du säker på att du vill radera gruppen?
hub.AssociateAGravatar=Koppla en <a href="http://www.gravatar.com" target="blank">Gravatar</a> till din e-postadress
hub.Availability=Tillgänglighet
hub.Block=Blockera
hub.Browse=Bläddra
hub.BrowseUsers=Bläddra i användarlistan
hub.Cancel=Avbryt
hub.CancelUpload=Avbryt uppladdningen
hub.CharactersLeft=bokstäver kvar
hub.ChooseALanguage=Välj ett språk
hub.Content=Innehåll
hub.CouldNotAddUser=Kunde inte lägga till användaren {0} till gruppen {0}
hub.CouldNotFindGroup=Kunde inte hitta någon grupp med id {0}
hub.CouldNotFindOrganization=Kunde inte hitta organisationen {0}
hub.CouldNotFindUser=Kunde inte hitta användaren {0}
hub.CouldNotRemoveDataset=Kunde inte ta bort Datasetet med id {0} från gruppen {0}
hub.CouldNotRemoveUser=Kunde inte ta bort användaren {0} från gruppen {0}
hub.CouldNotSaveGroup=Kunde inte spara gruppen, försök igen
hub.Create=Skapa
hub.CreateGroup=Skapa grupp
hub.Delete=Radera
hub.DeleteFiles=Radera filer
hub.Disable=Inaktivera
hub.Download=Ladda ner
hub.Edit=Redigera
hub.EditYourProfile=Redigera din profil
hub.Email=E-post
hub.EnlargeImage=Förstora bilden
hub.EnterANewPasswordBelow=Ange ett nytt lösenord nedan
hub.EnterASearchTerm=Skriv ett sökord och tryck [ENTER]
hub.EnterTheCodeYouSeeHere=Skriv in koden du ser här
hub.Error=Fel
hub.ErrorActivatingYourAccount.=Kunde inte aktivera ditt konto.
hub.ErrorChangingYourPassword=Kunde inte ändra ditt lösenord. Försök återställa det igen.
hub.ErrorCreatingYourAccount=Kunde inte skapa ditt konto, försök igen. Felmeddelande: {0}
hub.ErrorRemovingFile=Kunde inte ta bort filen,  Error removing file, ogiltigt id {0}
hub.ErrorResettingYourPassword=Kunde inte återställa ditt lösenord: {0}
hub.ErrorSavingTheme=Kunde inte spara tema {0}
hub.ErrorSavingYourProfile=Kunde inte spara din profil, försök igen
hub.First=Första
hub.FirstName=Förnamn
hub.FullName=Fullständigt namn
hub.FunFact=Roligt faktum
hub.GoTo=Gå till
hub.GroupList=Grupplista
hub.Hello=Hej
hub.Hi=Hej
hub.Home=Hem
hub.IForgotMyPassword=Jag har glömt mitt lösenord
hub.Identifier=Identifierare
hub.IfYouHaveForgottenYourPassword=Om du har glömt ditt lösenord kan du återställa det genom att skriva din e-postadress nedan
hub.Import=Importera
hub.InvalidCode=Ogiltig kod, skriv den igen
hub.Language=Språk
hub.Last=Sista
hub.LastName=Efternamn
hub.LaunchTheSIPCreatorBy=Starta SIP-Creator genom att klicka på logotypen till vänster. Din webbläsare kommer att vilja öppna en programfil som heter <strong>sip-creator.jnlp</strong> som kommer installeras på din dator. Du måste ha <strong>Java</strong> installerat på din dator. Varje gång du startar SIP-Creator kontrollerar den om det finns uppdateringar och uppdaterar automatiskt.
hub.Less=Mindre Less
hub.List=Lista
hub.ListAll=Lista allt
hub.ListOfHeritageObjects=Lista över kulturarvsobjekt
hub.ListOfHeritageObjectsFor=Lista över kulturarvsobjekt för {0}
hub.ListOfUsers=Lista över användare
hub.Load=Ladda
hub.Location=Placering
hub.LoggedInAs=Inloggad som
hub.Login=Logga in
hub.LoginIncorrect=Felaktig inloggning
hub.Logout=Logga ut
hub.LostPassword=Glömt lösenord
hub.Member=Medlem
hub.Members=Medlemmar
hub.More=Mer
hub.New=Ny
hub.Next=Nästa
hub.No=Nej
hub.NoAccountCouldBeFound=Inget konto kunde hittas med denna e-postadress
hub.NoProfileWasFound=Ingen profil hittades för användaren {0}
hub.NotAValidURL=Inte en giltig webbadress
hub.NotPublic=Ej publik
hub.NumberMembers={0} medlem/medlemmar
hub.NumberOfItems=Antal artiklar
hub.Options=Alternativ
hub.OrganizationAdministration=Organisations administrering
hub.OrganizationInformation=Organisations information
hub.Overview=Översikt
hub.Password=Lösenord
hub.PasswordIsRequired=Lösenord krävs
hub.PasswordsAreNotTheSame=Lösenorden är inte lika
hub.Phone=Telefon
hub.Place=Plats
hub.Places=Platser
hub.PoweredByDelving=Powered by DELVING.EU
hub.Preview=Förhandsgranska
hub.Previous=Föregående
hub.PreviousVersions=Tidigare versioner
hub.Print=Skriv ut
hub.Private=Privat
hub.ProfileActiveSince=Aktiv sedan
hub.ProfilePageFor=Profilsida för
hub.ProfileVisibleForNonconnectedUsers=Om du markerar det här alternativet, är din profil synlig för icke-anslutna användare
hub.Public=Publik
hub.Register=Registrera
hub.RegisterFor=Registrera för {0}
hub.RememberMe=Kom ihåg mig
hub.Remove=Ta bort
hub.RemovingAMemberWillAlso=Om du tar bort en medlem kommer den också att tas bort från alla grupper den är medlem i. Är du säker på att du vill fortsätta?
hub.RepeatPassword=Lösenord (repetera)
hub.Required=krävs
hub.Reset=Återställ
hub.ResetPassword=Återställ lösenord
hub.ResetPasswordTokenNotFound=Nyckeln för att återställa lösenordet hittades inte
hub.ReturnToResults=Återgå till resultatet
hub.SIPCreator=SIP-Creator
hub.Save=Spara
hub.SaveGroup=Spara grupp
hub.SaveProfile=Spara profil
hub.Scope=Omfattning
hub.Search=Sök
hub.SelectACollection=Välj en samling
hub.Share=Dela
hub.SorryNothingFound=Det verkar som det inte finns något att hitta just nu.
hub.StartUpload=Starta uppladdning
hub.State=Tillstånd
hub.Status=Status
hub.TheItemCannotBeDisplayed=Artikeln kan inte visas - {0}
hub.TheSIPCreatorIs=SIP-Creator är ett fristående verktyg som du kan använda för att hantera dina dataset. Det har funktioner som gör att du kan mappa alla befintliga XML-format till andra datadefinitioner som valts som mål för varje dataset individuellt. När datat är mappat och validerat, laddar SIP-Creator upp källdatat och mappningsfilen till Delving Culture Hub, så att mappningen kan göras där.
hub.Theme=Sidtema
hub.ThemeWithIdWasNotFound=Temat med id {0} kunde inte hittas
hub.ThereAreCurrentlyNoUsers=Det finns för närvarande inga användare i systemet (hur kom du in?)
hub.ThereIsAlreadyAUserWithThisEmailAddress=Det finns redan en användare med denna e-postadress
hub.ThereIsAlreadyAUserWithThisUsername=Det finns redan en användare med detta användarnamn
hub.ThisAccountIsNotActiveYet=Detta konto är inte aktiverat än. Aktivera kontot med hjälp av länken i registreringsmailet
hub.ThisObjectIsVisibleOnlyToYou=Detta objekt är bara synligt för dig. Om du vill att andra ska kunna söka och se det, kan du ändra objektets <a href="{0}"><strong>synlighets status</strong></a> till "Publik".
hub.ThisUsernameIsNotValid=Användarnamnet är inte giltig. Ett användarnamn kan endast innehålla små bokstäver, siffror och måste vara mellan 3 och 15 tecken långt.
hub.TypeHereToNarrowDown=Skriv här för att begränsa listan
hub.TypeHereToNarrowDownHelp=Skriv in ett värde för att filtrera listan. Tryck 'Spara' för att spara filtret. Tryck 'Återställ' för att ta bort filtret.
hub.Unlock=Lås upp
hub.User=Användare {0}
hub.UserWasNotFound=Användare {0} hittades inte
hub.Username=Användarnamn
hub.UsernameIsRequired=Användarnamn krävs
hub.ValueOutOfRange=Värdet är utanför godkänt intervall
hub.Visibility=Synlighet
hub.WarningOutdatedBrowser=<strong>Varning!</strong> Du har en föråldrad webbläsare. Denna webbplats kräver en modern, standard-kompatibel webbläsare för att fungera korrekt. Äldre webbläsare följer inte moderna standarderna och är också en allvarlig säkerhetsrisk för <em>din</em> dator.
hub.Website=Webbsida
hub.Welcome=Välkommen
hub.What=vad
hub.When=när
hub.Where=var
hub.Who=vem
hub.WithDigitalObject=Med digitalt objekt
hub.WithFullAccess=med full tillgång till allt
hub.WithRightsToModify=med rättigheter att ändra
hub.WithRightsToView=med rättigheter att visa
hub.WithoutDigitalObject=Utan digitalt objekt
hub.Yes=Ja
hub.YouDoNotHaveAccess=Vi ber om ursäkt, men du har inte behörighet hit
hub.YouWereLoggedOutSuccessfully=Du är nu utloggad
hub.YourAccountIsNotYetActive=Ditt konto är inte aktiverat än. Aktivera kontot med hjälp av länken i registreringsmailet
hub.YourAccountIsNowActive=Ditt konto är nu aktivt!
hub.YourAccountWasCreated=Ditt konto är nu skapat! Ett mail är skickat till {0} för aktivering
hub.YourBrowserNeedsToSupportCookies=Din webbläsare måste stödja cookies för att webbplatsen ska fungera korrekt.
hub.YourLinkedIn=Ditt linkedIn profilnamn, t ex johndoe
hub.YourPasswordHasBeenChanged=Ditt lösenord är nu ändrat
hub.YourPhoneNumber=Ditt telefonnummer
hub.YourProfile=Din profil
hub.YourTwitter=Ditt twitter användarnamn, t ex #johndoe
hubCompute=Beräkna
hubb.ALabelIs=En etikett är ett stycke text som du kan bifoga till ett objekt. En "fritext" etikett kan vara en beskrivande term. En "platsnamn" etikett bör avse en geografisk plats.
hubb.Action=Åtgärd
hubb.Actions=Åtgärder
hubb.AddComment=Lägg till kommentar
hubb.AddLabel=Lägg till etikett
hubb.Address=Adress
hubb.Administrator=Administratör
hubb.Administrators=Administratörer
hubb.AreYouSure=Är du säker?
hubb.AreYouSureYouWantToDelete=Är du säker på att du vill radera detta objekt?
hubb.Browse=Bläddra bland {0}
hubb.BrowseOf=Bläddra bland {0} av
hubb.BrowseOwnedBy=Bläddra bland {0} tillhörande
hubb.CancelUpload=Avbryt uppladdning
hubb.ChooseFile=Välj fil
hubb.City=Stad
hubb.Collaborators=Medarbetare
hubb.Collection=Samling
hubb.Collections=Samlingar
hubb.Comment=Kommentar
hubb.Comments=Kommentarer
hubb.Contact=Kontakt
hubb.ContactEmail=Kontakt e-post
hubb.ContactName=Kontakt namn
hubb.Content=Innehåll
hubb.CreateANew=Skapa en ny {0}
hubb.CreatingACaptivatingNarrative=Skapa en fängslande berättelse är ibland det enda sättet att ge kulturföremål sammanhanget de förtjänar. Ofta gör deras beskrivningar dem inte rättvisa, men att använda dem i en berättelse med några av dina kulturskatter skulle kanske kunna skapa något mycket bättre. Denna webbplats gör det lättare för oss att bygga dessa berättelser och göra dem tillgängliga för alla att ta del av.
hubb.Creator=Skapare
hubb.DateCreated=Skapad datum
hubb.DateModified=Ändrad datum
hubb.Description=Beskrivning
hubb.Email=E-post
hubb.EndYear=Slut år
hubb.Fax=Fax
hubb.FileName=Filnamn
hubb.FileSize=Filstorlek
hubb.FreeTextLabel=Fritext etikett
hubb.GeographicalArea=Geografiskt område
hubb.Group=Grupp
hubb.Groups=Grupper
hubb.HeritageObject=Kulturarvsobjekt
hubb.ImageDocumentUpload=Bild/dokument uppladdning
hubb.Instant=Omedelbar
hubb.Keyword=Nyckelord
hubb.Keywords=Nyckelord
hubb.Label=Etikett
hubb.Labels=Etiketter
hubb.LandingPage=Målsida
hubb.Measurements=Mått
hubb.MissionStatement=verksamhetsidé
hubb.Municipality=Kommun
hubb.Museum=Museum
hubb.Museums=Museum
hubb.Name=Namn
hubb.Object=Objekt
hubb.Objects.heritage=Kulturarvsobjekt
hubb.Objects=Objekt
hubb.Organization=Organisation
hubb.Organizations=Organisationer
hubb.Owner=Ägare
hubb.Place=Plats
hubb.PlaceNameLabel=Platsnamn etikett
hubb.PostalCode=Postnummer
hubb.Provider=Leverantör
hubb.Province=Region
hubb.RelatedItems=Relaterade objekt
hubb.Resources=Resurser
hubb.SitePage=Webbsida
hubb.SitePages=Webbsidor
hubb.StartUpload=Starta uppladdning
hubb.StartYear=Start år
hubb.Stories=Historier
hubb.Story=Historia
hubb.ThereAreCurrentlyNoAvailable=Det finns för tillfället ingen {0} tillgänglig
hubb.ThereIsCurrentlyNoAvailable=Det finns för tillfället ingen {0} tillgänglig
hubb.ThisGroupGrants=Denna grupp beviljar
hubb.Thumbnail=Tumnagel
hubb.Title=Titel
hubb.URL=URL
hubb.UploadedFiles=Uppladdade filer
hubb.User=Användare
hubb.Users=Användare
hubb.Version=Version
hubnode.ANodeWithTheSameNodeIdentifier=En nod med samma nod id finns redan
hubnode.AreYouSureYouWantToDeleteThisHubNode=Är du säker på att du vill radera denna virtuella nod och data kopplat till den?
hubnode.CreateHubNode=Skapa Hub nod
hubnode.HubNode=Hub nod
hubnode.HubNodes=Hub noder
hubnode.InvalidNodeName=Ogiltigt nodnamn: kan bara innehålla bokstäver och mellanslag
hubnode.ListHubNodes=Lista över Hub noder
hubnode.NodeIdentifier=Nod id
hubnode.NodeName=Nodnamn
hubnode.OrganizationIdentifier=Organisations id
hubnode.ThisOrganizationDoesntExist=Denna organisation finns inte inlagd. Kontakta support@delving.eu för hjälp.
lang.Dutch=Holländska (nl)
lang.English=Engelska (en)
lang.Norwegian=Norska (no)
lang.NorwegianBokmal=Norska bokmål (nb)
mail.InOrderToResetYourPassword=För att återställa ditt lösenord för {0}, tryck på länken nedan
mail.YourAccountHasBeenBlocked=Ditt konto har blockerats på grund av att det innehåll du har skrivit in inte bedöms vara lämplig för den här webbplatsen. Om du tycker detta är fel, kontakta {0}.
mail.YourAccountHasBeenBlockedSubject=Ditt konto har blockerats
mail.YourAccountHasBeenCreated=Ditt konto för {0} har skapats. För att aktivera ditt konto, klicka på länken nedan
metadata.abm.aboutPerson=Om personen
metadata.abm.address=Adress
metadata.abm.contentProvider=Innehålls leverantör
metadata.abm.county=Län
metadata.abm.dataProvider=Dataleverantör
metadata.abm.digitised=Digitaliserad
metadata.abm.geo=Geo-koordinater
metadata.abm.landedProperty=Fast egendom
metadata.abm.latitude=Latitud
metadata.abm.longitude=Longitud
metadata.abm.municipality=Kommun
metadata.abm.namedPlace=Platsnamn
metadata.coll.AATCategories=AAT kategorier
metadata.coll.Administrators=Administratörer
metadata.coll.Borrowed=Lånad
metadata.coll.EarliestWorkFromCollection=Tidigaste verk från samlingen
metadata.coll.FromCoreCollection=Från huvudsamling
metadata.coll.GeographicalRelevance=Geografisk relevans
metadata.coll.MostRecentWorkFromCollection=Det senaste verket från samlingen
metadata.coll.Museum=Museum
metadata.coll.NumberOfObjects=Antal objekt
metadata.coll.RelationToCoreCollection=Relation till huvudsamling
metadata.coll.Strength=Styrka
metadata.coll.Total=Total
metadata.dc.contributor=Givare
metadata.dc.coverage=Täckning
metadata.dc.creator=Skapare
metadata.dc.date=Datum
metadata.dc.description=Beskrivning
metadata.dc.format=Format
metadata.dc.identifier=Identifierare
metadata.dc.language=Språk
metadata.dc.publisher=Utgivare
metadata.dc.relation=Relation
metadata.dc.rights=Rättigheter
metadata.dc.source=Källa
metadata.dc.subject=Ämne
metadata.dc.title=Titel
metadata.dc.type=Typ
metadata.dcterms.alternative=Alternativ Titel
metadata.dcterms.conformsTo=Uppfyller
metadata.dcterms.created=Datum skapad
metadata.dcterms.extent=Omfattning
metadata.dcterms.hasFormat=Har format
metadata.dcterms.hasPart=Har del
metadata.dcterms.hasVersion=Har version
metadata.dcterms.isFormatOf=Är av formatet
metadata.dcterms.isPartOf=Är del av
metadata.dcterms.isReferencedBy=Refereras av
metadata.dcterms.isReplacedBy=Ersätts av
metadata.dcterms.medium=Medium
metadata.dcterms.provenance=Proveniens
metadata.dcterms.references=Referenser
metadata.dcterms.replaces=Ersätts
metadata.dcterms.requires=Kräver
metadata.dcterms.rightsHolder=Rättighetsinnehavare
metadata.dcterms.spatialCoverage=Geografisk täckning
metadata.dcterms.temporalCoverage=Tidsmässig täckning
metadata.delving.collection=Samling
metadata.delving.creator=Skapad av
metadata.delving.description=Beskrivning
metadata.delving.dimensions=Dimensioner
metadata.delving.fullTextObjectUrl=Fulltext
metadata.delving.hasDigitalObject=Har bild
metadata.delving.owner=Dataägare
metadata.delving.provider=Dataleverantör
metadata.delving.recordType=Objekttyp
metadata.delving.title=Titel
metadata.europeana.collectionName=Samlingsnamn
metadata.europeana.collectionTitle=Samlingstitel
metadata.europeana.country=Land
metadata.europeana.dataProvider=Dataleverantör
metadata.europeana.isShownAt=Extern målsida
metadata.europeana.isShownBy=Extern url till det digitala objektet
metadata.europeana.language=Språk
metadata.europeana.object=Objekt
metadata.europeana.provider=Leverantör
metadata.europeana.rights=Rättigheter
metadata.europeana.type=Typ
metadata.europeana.uri=Europeana URI
metadata.europeana.year=År
metadata.icn.acceptedStateCharges=Godkända statliga avgifter
metadata.icn.acceptedStateChargesReason=Anledning till vedertagna statliga avgifter
metadata.icn.acquiredWithHelpFrom=Förvärvad med hjälp av
metadata.icn.acquisitionMeans=Mening med förvärv
metadata.icn.acquisitionYear=Förvärvat år
metadata.icn.collection=Samling
metadata.icn.collectionPart=Del
metadata.icn.collectionType=Samlingstyp
metadata.icn.creatorYearOfBirth=Skapare född
metadata.icn.creatorYearOfDeath=Skapare död
metadata.icn.currentLocation=Nuvarande placering
metadata.icn.expulsionMeans=Mening med uteslutning
metadata.icn.expulsionYear=Utesluten år
metadata.icn.legalStatus=Rättslig status
metadata.icn.location=Placering
metadata.icn.material=Material
metadata.icn.physicalState=Fysiskt tillstånd
metadata.icn.previousLocation=Tidigare placering
metadata.icn.province=Region
metadata.icn.purchasePrice=Inköpspris
metadata.icn.technique=Teknik
metadata.lido.actorInRole=Aktör i händelsen
metadata.lido.actor.roleActor=Roll
metadata.lido.administrativeMetadata.recordWrap=Objekt
metadata.lido.administrativeMetadata.recordWrap.recordID=ObjektId
metadata.lido.administrativeMetadata.resourceWrap=Resurs
metadata.lido.administrativeMetadata.rightsWorkWrap=Rättigheter
metadata.lido.category=Kategori
metadata.lido.conceptID=KonceptId
metadata.lido.displayDate=Datum
metadata.lido.displaySubject=Ämne
metadata.lido.displayPlace=Plats
metadata.lido.earliestDate=Tidigaste datum
metadata.lido.eventType=Typ av händelse
metadata.lido.eventWrap=Händelser
metadata.lido.event.eventActor=Aktör
metadata.lido.genderActor=Kön
metadata.lido.latestDate=Senaste datum
metadata.lido.legalBodyName=Juridiskt namn
metadata.lido.legalBodyWeblink=Juridisk person webbplats
metadata.lido.lidoRecId=PostId
metadata.lido.lidoRecId.source=Källa
metadata.lido.nationalityActor.term=Nationalitet
metadata.lido.objectClassificationWrap=Klassificering
metadata.lido.objectIdentificationWrap=Identitetsnummer
metadata.lido.objectRelationWrap.subjectWrap=Ämnen
metadata.lido.recordInfoID=URI
metadata.lido.recordInfoLink=Webbsida
metadata.lido.recordType=Objekttyp
metadata.lido.resourceType=Resurstyp
metadata.lido.rightsType=Typ av rättighet
metadata.lido.subject.subjectConcept.term=Term
metadata.lido.titleSet=Titel
metadata.lido.type=Typ
metadata.lido.workID=VerkId
metadata.text=Text
metadata.tib.citName=CIT samlingsnamn
metadata.tib.citOldId=CIT post id
metadata.tib.collection=Samling
metadata.tib.collectionPart=Under-samling
metadata.tib.color=färg
metadata.tib.creatorBirthYear=Födelseår
metadata.tib.creatorDeathYear=Dödsår
metadata.tib.creatorRole=Skapare roll
metadata.tib.date=Datum
metadata.tib.deepZoomUrl=URL för DeepZoom bild
metadata.tib.design=Design
metadata.tib.dimension=Dimension
metadata.tib.event=Händelse
metadata.tib.exhibition=Utställning
metadata.tib.formatted=Formaterad
metadata.tib.fullTextObjectUrl=URL till full-text sökbara objekt
metadata.tib.location=Geo-placering
metadata.tib.material=Material
metadata.tib.objectNumber=Inventarienummer
metadata.tib.objectSoort=Objekttyp
metadata.tib.pageEnd=Sista sidan
metadata.tib.pageStart=Startsidan
metadata.tib.pages=Sidor
metadata.tib.period=Period
metadata.tib.person=Person
metadata.tib.place=Plats
metadata.tib.productionEnd=Produktion slutdatum
metadata.tib.productionPeriod=Produktion period
metadata.tib.productionStart=Produktion startdatum
metadata.tib.region=Region
metadata.tib.subjectDepicted=Avbildat ämne
metadata.tib.technique=Teknik
metadata.tib.theme=Tema
metadata.tib.thumbLarge=Stor tumnagel
metadata.tib.thumbSmall=Liten tumnagel
metadata.tib.vindplaats=Fysisk placering
metadata.tib.year=År
metadata.type.All=Alla
metadata.type.Images=Bilder
metadata.type.Sounds=Ljud
metadata.type.Texts=Texter
metadata.type.Video=Video
metadata.type.Videos=Videor
mediator.Mediator=Förmedlare
sdu.AreYouSureYouWantToDelete=Är du säker på att du vill radera detta objekt?
sdu.DocumentUpload=Dokument uppladdning
sdu.ListOfUploadedDocuments=Lista på uppladdade dokument
sdu.UploadDocument=Ladda upp dokument
search.CannotConnectToTheSearchBackend=Kan inte ansluta till sökmotorn
search.Collection=Samling
search.Facets=Fasetter
search.FoundResults=Hittade {0} poster
search.ObjectType=Objekt typ
search.Provider=Leverantör
search.QueryIsNotValid=Sökning på "{0}" är inte giltig. Försök igen.
search.RefineYourSearch=Förfina din sökning
search.ResultsFor=Sökresultat för
search.ResultsOf=Resultat <strong>{0} - {1}</strong> av <strong>{2}</strong>
search.SortBy=Sortera på
search.ViewInOriginalContext=Visa i original kontext
search.Year=År
stats.History=Historia
stats.NumberOfRecords=Antal poster
stats.Statistics=Statistik
stats.WithGeographicalData=Med geografiskt data
stats.WithLandingPages=Med målsida
stats.WithObjects=Med objekt
stats.WithoutObjects=Utan objekt
